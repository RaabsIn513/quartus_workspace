library verilog;
use verilog.vl_types.all;
entity blockEd is
    port(
        pin_name1       : out    vl_logic;
        Input_sw        : in     vl_logic
    );
end blockEd;
