library verilog;
use verilog.vl_types.all;
entity ALU_TestBench is
end ALU_TestBench;
