
// Implements a simple Nios II system for the DE-series board.
// Inputs: SW7¡0 are parallel port inputs to the Nios II system
// CLOCK_50 is the system clock
// KEY0 is the active-low system reset
// Outputs: LEDG7¡0 are parallel port outputs from the Nios II system
module de0_tutorial (SW, KEY, CLOCK_50, LEDG);
input [7:0] SW;
input [0:0] KEY;
input CLOCK_50;
output [7:0] LEDG;
// Instantiate the Nios II system module generated by the SOPC Builder:
// nios_system (clk_0, reset_n, out_port_from_the_LEDs, in_port_to_the_Switches)
nios_system NiosII (CLOCK_50, KEY[0], LEDG, SW);

endmodule
