library verilog;
use verilog.vl_types.all;
entity usePC_TestBench is
end usePC_TestBench;
