library verilog;
use verilog.vl_types.all;
entity aTestBench is
end aTestBench;
