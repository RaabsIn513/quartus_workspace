library verilog;
use verilog.vl_types.all;
entity PC_TestBench is
end PC_TestBench;
