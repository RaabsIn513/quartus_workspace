library verilog;
use verilog.vl_types.all;
entity Memory_TestBench is
end Memory_TestBench;
