library verilog;
use verilog.vl_types.all;
entity TOP_TestBench is
end TOP_TestBench;
