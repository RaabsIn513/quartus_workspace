library verilog;
use verilog.vl_types.all;
entity clkDiv_TestBench is
end clkDiv_TestBench;
