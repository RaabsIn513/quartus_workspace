library verilog;
use verilog.vl_types.all;
entity Adder_TestBench is
end Adder_TestBench;
