library verilog;
use verilog.vl_types.all;
entity aTB is
end aTB;
