library verilog;
use verilog.vl_types.all;
entity blockEd is
    port(
        in_pin          : in     vl_logic;
        out_pin         : out    vl_logic
    );
end blockEd;
