library verilog;
use verilog.vl_types.all;
entity cpu_0_nios2_performance_monitors is
end cpu_0_nios2_performance_monitors;
