module proc_TestBench;
  //proc( clk, reset, LCD, lcdRS, lcdRW, lcdEn, LED );
  
  reg clock, rst;
  wire[7:0] LCD;
  wire lcdRW, lcdEn, LEDtb, lcdRS;
  
  initial begin
    #2 clock <= 1'b0;
    #10 rst <= 1'b0;
    #20 rst <= 1'b1;
  end
  
  always begin
    #5 clock <= !clock;
  end
  //proc( clk, reset, LCD, lcdRS, lcdRW, lcdEn, LED );
  proc U0( clock, rst, LCD, lcdRS, lcdRW, lcdEn, LEDtb );

  
endmodule