library verilog;
use verilog.vl_types.all;
entity useClkDive_TestBench is
end useClkDive_TestBench;
