library verilog;
use verilog.vl_types.all;
entity LCD_Driver_TestBench is
end LCD_Driver_TestBench;
