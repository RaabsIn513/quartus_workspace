library verilog;
use verilog.vl_types.all;
entity proc_TestBench is
end proc_TestBench;
