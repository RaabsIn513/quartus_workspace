library verilog;
use verilog.vl_types.all;
entity ALU_testBench is
end ALU_testBench;
