library verilog;
use verilog.vl_types.all;
entity cpu_0_data_master_arbitrator is
    port(
        Switches_s1_readdata_from_sa: in     vl_logic_vector(31 downto 0);
        clk             : in     vl_logic;
        clocks_0_avalon_clocks_slave_readdata_from_sa: in     vl_logic_vector(7 downto 0);
        cpu_0_data_master_address: in     vl_logic_vector(24 downto 0);
        cpu_0_data_master_byteenable_sdram_0_s1: in     vl_logic_vector(1 downto 0);
        cpu_0_data_master_granted_Switches_s1: in     vl_logic;
        cpu_0_data_master_granted_clocks_0_avalon_clocks_slave: in     vl_logic;
        cpu_0_data_master_granted_cpu_0_jtag_debug_module: in     vl_logic;
        cpu_0_data_master_granted_greenLEDS_s1: in     vl_logic;
        cpu_0_data_master_granted_jtag_uart_0_avalon_jtag_slave: in     vl_logic;
        cpu_0_data_master_granted_onchip_memory2_0_s1: in     vl_logic;
        cpu_0_data_master_granted_sdram_0_s1: in     vl_logic;
        cpu_0_data_master_granted_timer_0_s1: in     vl_logic;
        cpu_0_data_master_qualified_request_Switches_s1: in     vl_logic;
        cpu_0_data_master_qualified_request_clocks_0_avalon_clocks_slave: in     vl_logic;
        cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module: in     vl_logic;
        cpu_0_data_master_qualified_request_greenLEDS_s1: in     vl_logic;
        cpu_0_data_master_qualified_request_jtag_uart_0_avalon_jtag_slave: in     vl_logic;
        cpu_0_data_master_qualified_request_onchip_memory2_0_s1: in     vl_logic;
        cpu_0_data_master_qualified_request_sdram_0_s1: in     vl_logic;
        cpu_0_data_master_qualified_request_timer_0_s1: in     vl_logic;
        cpu_0_data_master_read: in     vl_logic;
        cpu_0_data_master_read_data_valid_Switches_s1: in     vl_logic;
        cpu_0_data_master_read_data_valid_clocks_0_avalon_clocks_slave: in     vl_logic;
        cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module: in     vl_logic;
        cpu_0_data_master_read_data_valid_greenLEDS_s1: in     vl_logic;
        cpu_0_data_master_read_data_valid_jtag_uart_0_avalon_jtag_slave: in     vl_logic;
        cpu_0_data_master_read_data_valid_onchip_memory2_0_s1: in     vl_logic;
        cpu_0_data_master_read_data_valid_sdram_0_s1: in     vl_logic;
        cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register: in     vl_logic;
        cpu_0_data_master_read_data_valid_timer_0_s1: in     vl_logic;
        cpu_0_data_master_requests_Switches_s1: in     vl_logic;
        cpu_0_data_master_requests_clocks_0_avalon_clocks_slave: in     vl_logic;
        cpu_0_data_master_requests_cpu_0_jtag_debug_module: in     vl_logic;
        cpu_0_data_master_requests_greenLEDS_s1: in     vl_logic;
        cpu_0_data_master_requests_jtag_uart_0_avalon_jtag_slave: in     vl_logic;
        cpu_0_data_master_requests_onchip_memory2_0_s1: in     vl_logic;
        cpu_0_data_master_requests_sdram_0_s1: in     vl_logic;
        cpu_0_data_master_requests_timer_0_s1: in     vl_logic;
        cpu_0_data_master_write: in     vl_logic;
        cpu_0_data_master_writedata: in     vl_logic_vector(31 downto 0);
        cpu_0_jtag_debug_module_readdata_from_sa: in     vl_logic_vector(31 downto 0);
        d1_Switches_s1_end_xfer: in     vl_logic;
        d1_clocks_0_avalon_clocks_slave_end_xfer: in     vl_logic;
        d1_cpu_0_jtag_debug_module_end_xfer: in     vl_logic;
        d1_greenLEDS_s1_end_xfer: in     vl_logic;
        d1_jtag_uart_0_avalon_jtag_slave_end_xfer: in     vl_logic;
        d1_onchip_memory2_0_s1_end_xfer: in     vl_logic;
        d1_sdram_0_s1_end_xfer: in     vl_logic;
        d1_timer_0_s1_end_xfer: in     vl_logic;
        greenLEDS_s1_readdata_from_sa: in     vl_logic_vector(31 downto 0);
        jtag_uart_0_avalon_jtag_slave_irq_from_sa: in     vl_logic;
        jtag_uart_0_avalon_jtag_slave_readdata_from_sa: in     vl_logic_vector(31 downto 0);
        jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa: in     vl_logic;
        onchip_memory2_0_s1_readdata_from_sa: in     vl_logic_vector(31 downto 0);
        registered_cpu_0_data_master_read_data_valid_clocks_0_avalon_clocks_slave: in     vl_logic;
        registered_cpu_0_data_master_read_data_valid_onchip_memory2_0_s1: in     vl_logic;
        reset_n         : in     vl_logic;
        sdram_0_s1_readdata_from_sa: in     vl_logic_vector(15 downto 0);
        sdram_0_s1_waitrequest_from_sa: in     vl_logic;
        timer_0_s1_irq_from_sa: in     vl_logic;
        timer_0_s1_readdata_from_sa: in     vl_logic_vector(15 downto 0);
        cpu_0_data_master_address_to_slave: out    vl_logic_vector(24 downto 0);
        cpu_0_data_master_dbs_address: out    vl_logic_vector(1 downto 0);
        cpu_0_data_master_dbs_write_16: out    vl_logic_vector(15 downto 0);
        cpu_0_data_master_irq: out    vl_logic_vector(31 downto 0);
        cpu_0_data_master_no_byte_enables_and_last_term: out    vl_logic;
        cpu_0_data_master_readdata: out    vl_logic_vector(31 downto 0);
        cpu_0_data_master_waitrequest: out    vl_logic
    );
end cpu_0_data_master_arbitrator;
