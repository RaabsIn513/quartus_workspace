library verilog;
use verilog.vl_types.all;
entity LCD_TestBench is
end LCD_TestBench;
